`include "sv/apb_master_driver_orig.sv"
